//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel,
  output [3:0] y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

  // Task:
  // Implement mux_4_1 using three instances of mux_2_1

  logic [3:0] d32, d10;

  mux_2_1 i0_mux (
    .d1  ( d3      ),
    .d0  ( d2      ),
    .sel ( sel [0] ),
    .y   ( d32     )
  );

  mux_2_1 i1_mux (
    .d1  ( d1      ),
    .d0  ( d0      ),
    .sel ( sel [0] ),
    .y   ( d10     )
  );

  mux_2_1 i2_mux (
    .d1  ( d32     ),
    .d0  ( d10     ),
    .sel ( sel [1] ),
    .y   ( y       )
  );

endmodule
